/*
+ Project   : Emulator Graduation Project 2018 ASU-CSE
+ Module    : Weight ROM
+ Abstract  : The ROM storing the weights of a single neuron
+ Notes     : 
  - Each ALU has its own ROM that stores the its corresponding weights of a specific neuron
  - The address counter reset is sync. with the clock edge
  - The memory .TXT file should store the weigh values IN BINARY REPRESENTATION
  - The memory is single ported and read only; with an internal address pointer that auto increments each cycle
  - Loading the memory is done by specifying the external text file generated by the pre-processor containing
    the weights of one neuron
  - The FILE_NAME content must have a total number of bits / word = BIT_WIDTH+EXTRA_BITS
*/

`ifndef WEIGHTS_ROM_
`define WEIGHTS_ROM_
`default_nettype none
`include "definitions.v"

module WEIGHTS_ROM #(
  parameter BIT_WIDTH = 32,               // The floating point size in bits
  parameter EXTRA_BITS = 2,               // Flopoco Floating point extra two bits. CAN ONLY have the values [0 OR 2]
  parameter DEPTH =  4,                   // Memory depth [Number of elements or words in memory]
  parameter MEM_DIR = `MEM_DIR,           // Directory holding all memory files
  parameter PTR_RESET_BASE = 0,           // Counter reset value
  parameter FILE_NAME = "init.txt"    // The .txt file holding the weights to be stored into the memory IN BINARY REPRESENTATION
)
(
  input wire                                CLK,        // Sync. clock
  input wire                                RESET,      // Resetting the address pointer back to zero [the first weight]
  output wire                               ACC_EN,     // ALU signal for enabling/disabling accumulator based on the current address
  output reg [BIT_WIDTH + EXTRA_BITS - 1:0] MEM_OUT     // The weight participating in the MACC operation
);

  // Internal wires, reg declaration area
  reg [BIT_WIDTH + EXTRA_BITS - 1:0] weight_memory [0:DEPTH-1];       // Memory holding all the neuron weights
  reg [$clog2(DEPTH)-1: 0] address_ptr;                               // Address pointer
  // Internal wires assignment
  assign ACC_EN = address_ptr!=1;
  
  // Memory filling routine
  /*ANY EXTRA SYNTHESIS FLAGS/COMMANDS SHOULD BE PLACED HERE */
  initial begin
    $readmemb(FILE_NAME, weight_memory);
  end

  // Functional blocks
  always @(posedge CLK ) begin
    if(RESET) begin
      address_ptr <= PTR_RESET_BASE;//0;
    end
    else begin
      if (address_ptr == (DEPTH-1)) begin
        address_ptr <=0;
      end
      else begin
        address_ptr <= address_ptr +1;
      end
    end
    MEM_OUT <= weight_memory[address_ptr];
  end

endmodule // WEIGHTS_ROM
`endif